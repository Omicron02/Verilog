module not1(b,a);
    input a;
    output b;
    assign b=~a;
endmodule 